`define KNN_ADDR_W 3  //address width
`define KNN_WDATA_W 1 //write data width
`ifndef DATA_W
 `define DATA_W 32      //cpu data width
`endif

`ifndef DATASET_SIZE
 `define DATASET_SIZE 100      //Dataset number (abitrario)
`endif
